module counter(

);